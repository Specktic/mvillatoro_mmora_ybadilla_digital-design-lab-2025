package OpCodeEnum;

	typedef enum {
		Add,
		Sub,
		Mult,
		Div,
		Mod,
		And,
		Or,
		Xor,
		LShift,
		RShift
	} OpCode;

endpackage