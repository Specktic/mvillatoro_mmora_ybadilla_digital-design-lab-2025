/*Testbench*/